`ifndef IMM_TYPE_MAC_H
`define IMM_TYPE_MAC_H

`define IMM_TYPE_I    3'b000
`define IMM_TYPE_S    3'b001
`define IMM_TYPE_B    3'b010
`define IMM_TYPE_U    3'b011
`define IMM_TYPE_J    3'b100
`define IMM_TYPE_NONE 3'b111

`endif
