`ifndef RV32I_LSU_I_MAC_H
`define RV32I_LSU_I_MAC_H

`define RV32I_LSU_I_OPCODE 7'b0000011

`define RV32I_LSU_I_F3_LB  3'h0
`define RV32I_LSU_I_F3_LH  3'h1
`define RV32I_LSU_I_F3_LW  3'h2
`define RV32I_LSU_I_F3_LBU 3'h4
`define RV32I_LSU_I_F3_LHU 3'h5

`endif
