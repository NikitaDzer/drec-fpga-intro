`ifndef ALU_A_SEL_MAC_H
`define ALU_A_SEL_MAC_H

`define ALU_A_SEL_REG 1'b0
`define ALU_A_SEL_IMM 1'b1

`endif
