`ifndef RV32I_ALU_I_MAC_H
`define RV32I_ALU_I_MAC_H

`define RV32I_ALU_I_OPCODE 7'b0010011

`define RV32I_ALU_I_F3_ADDI  3'h0
`define RV32I_ALU_I_F3_XORI  3'h4
`define RV32I_ALU_I_F3_ORI   3'h6
`define RV32I_ALU_I_F3_ANDI  3'h7
`define RV32I_ALU_I_F3_SLLI  3'h1
`define RV32I_ALU_I_F3_SRLI  3'h5
`define RV32I_ALU_I_F3_SRAI  3'h5
`define RV32I_ALU_I_F3_SLTI  3'h2
`define RV32I_ALU_I_F3_SLTIU 3'h3

`endif
