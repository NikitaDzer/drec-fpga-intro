`ifndef WB_SEL_MAC_H
`define WB_SEL_MAC_H

`define WB_SEL_ALU      2'b00
`define WB_SEL_LSU      2'b01
`define WB_SEL_PC32_INC 2'b10
`define WB_SEL_IMM      2'b11

`endif
