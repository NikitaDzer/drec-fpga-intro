module copy_bit (
    input  wire i_bit,
    output wire o_bit
);

assign o_bit = i_bit;

endmodule
