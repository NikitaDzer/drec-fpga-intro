`ifndef RV32I_CBU_J_MAC_H
`define RV32I_CBU_J_MAC_H

`define RV32I_CBU_J_OPCODE_JAL 7'b1101111

`endif
