`ifndef BU_MAC_H
`define BU_MAC_H

`define BU_BEQ  3'b000
`define BU_BNE  3'b001
`define BU_BLT  3'b010
`define BU_BGE  3'b011
`define BU_BLTU 3'b100
`define BU_BGEU 3'b101
`define BU_PT   3'b110
`define BU_NONE 3'b111

`endif
