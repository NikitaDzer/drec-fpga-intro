`ifndef RV32I_LSU_S_MAC_H
`define RV32I_LSU_S_MAC_H

`define RV32I_LSU_S_OPCODE 7'b0100011

`define RV32I_LSU_S_F3_SB 3'h0
`define RV32I_LSU_S_F3_SH 3'h1
`define RV32I_LSU_S_F3_SW 3'h2

`endif
