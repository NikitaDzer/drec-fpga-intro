`ifndef ALU_B_SEL_MAC_H
`define ALU_B_SEL_MAC_H

`define ALU_B_SEL_REG  2'b00
`define ALU_B_SEL_IMM  2'b01
`define ALU_B_SEL_PC32 2'b10

`endif
