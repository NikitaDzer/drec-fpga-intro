`ifndef RV32I_CBU_B_MAC_H
`define RV32I_CBU_B_MAC_H

`define RV32I_CBU_B_OPCODE 7'b1100011

`define RV32I_CBU_B_F3_BEQ  3'h0
`define RV32I_CBU_B_F3_BNE  3'h1
`define RV32I_CBU_B_F3_BLT  3'h4
`define RV32I_CBU_B_F3_BGE  3'h5
`define RV32I_CBU_B_F3_BLTU 3'h6
`define RV32I_CBU_B_F3_BGEU 3'h7

`endif
